// system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system (
		input  wire        reset_reset_n,    //      reset.reset_n
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		input  wire        sys_clk_clk       //    sys_clk.clk
	);

	wire         pll_0_outclk0_clk;                                           // pll_0:outclk_0 -> [SHA_0:clk, SHA_1:clk, SHA_2:clk, SHA_3:clk, SHA_4:clk, SHA_5:clk, SHA_6:clk, SHA_7:clk, SHA_8:clk, SHA_9:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, irq_synchronizer_004:receiver_clk, irq_synchronizer_005:receiver_clk, irq_synchronizer_006:receiver_clk, irq_synchronizer_007:receiver_clk, irq_synchronizer_008:receiver_clk, irq_synchronizer_009:receiver_clk, mm_interconnect_0:pll_0_outclk0_clk, rst_controller:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [26:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_sha_0_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_0_avalon_slave_0_chipselect -> SHA_0:cs
	wire  [31:0] mm_interconnect_0_sha_0_avalon_slave_0_readdata;             // SHA_0:read_data -> mm_interconnect_0:SHA_0_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_0_avalon_slave_0_address;              // mm_interconnect_0:SHA_0_avalon_slave_0_address -> SHA_0:address
	wire         mm_interconnect_0_sha_0_avalon_slave_0_write;                // mm_interconnect_0:SHA_0_avalon_slave_0_write -> SHA_0:we
	wire  [31:0] mm_interconnect_0_sha_0_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_0_avalon_slave_0_writedata -> SHA_0:write_data
	wire         mm_interconnect_0_sha_1_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_1_avalon_slave_0_chipselect -> SHA_1:cs
	wire  [31:0] mm_interconnect_0_sha_1_avalon_slave_0_readdata;             // SHA_1:read_data -> mm_interconnect_0:SHA_1_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_1_avalon_slave_0_address;              // mm_interconnect_0:SHA_1_avalon_slave_0_address -> SHA_1:address
	wire         mm_interconnect_0_sha_1_avalon_slave_0_write;                // mm_interconnect_0:SHA_1_avalon_slave_0_write -> SHA_1:we
	wire  [31:0] mm_interconnect_0_sha_1_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_1_avalon_slave_0_writedata -> SHA_1:write_data
	wire         mm_interconnect_0_sha_2_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_2_avalon_slave_0_chipselect -> SHA_2:cs
	wire  [31:0] mm_interconnect_0_sha_2_avalon_slave_0_readdata;             // SHA_2:read_data -> mm_interconnect_0:SHA_2_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_2_avalon_slave_0_address;              // mm_interconnect_0:SHA_2_avalon_slave_0_address -> SHA_2:address
	wire         mm_interconnect_0_sha_2_avalon_slave_0_write;                // mm_interconnect_0:SHA_2_avalon_slave_0_write -> SHA_2:we
	wire  [31:0] mm_interconnect_0_sha_2_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_2_avalon_slave_0_writedata -> SHA_2:write_data
	wire         mm_interconnect_0_sha_3_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_3_avalon_slave_0_chipselect -> SHA_3:cs
	wire  [31:0] mm_interconnect_0_sha_3_avalon_slave_0_readdata;             // SHA_3:read_data -> mm_interconnect_0:SHA_3_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_3_avalon_slave_0_address;              // mm_interconnect_0:SHA_3_avalon_slave_0_address -> SHA_3:address
	wire         mm_interconnect_0_sha_3_avalon_slave_0_write;                // mm_interconnect_0:SHA_3_avalon_slave_0_write -> SHA_3:we
	wire  [31:0] mm_interconnect_0_sha_3_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_3_avalon_slave_0_writedata -> SHA_3:write_data
	wire         mm_interconnect_0_sha_4_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_4_avalon_slave_0_chipselect -> SHA_4:cs
	wire  [31:0] mm_interconnect_0_sha_4_avalon_slave_0_readdata;             // SHA_4:read_data -> mm_interconnect_0:SHA_4_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_4_avalon_slave_0_address;              // mm_interconnect_0:SHA_4_avalon_slave_0_address -> SHA_4:address
	wire         mm_interconnect_0_sha_4_avalon_slave_0_write;                // mm_interconnect_0:SHA_4_avalon_slave_0_write -> SHA_4:we
	wire  [31:0] mm_interconnect_0_sha_4_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_4_avalon_slave_0_writedata -> SHA_4:write_data
	wire         mm_interconnect_0_sha_5_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_5_avalon_slave_0_chipselect -> SHA_5:cs
	wire  [31:0] mm_interconnect_0_sha_5_avalon_slave_0_readdata;             // SHA_5:read_data -> mm_interconnect_0:SHA_5_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_5_avalon_slave_0_address;              // mm_interconnect_0:SHA_5_avalon_slave_0_address -> SHA_5:address
	wire         mm_interconnect_0_sha_5_avalon_slave_0_write;                // mm_interconnect_0:SHA_5_avalon_slave_0_write -> SHA_5:we
	wire  [31:0] mm_interconnect_0_sha_5_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_5_avalon_slave_0_writedata -> SHA_5:write_data
	wire         mm_interconnect_0_sha_6_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_6_avalon_slave_0_chipselect -> SHA_6:cs
	wire  [31:0] mm_interconnect_0_sha_6_avalon_slave_0_readdata;             // SHA_6:read_data -> mm_interconnect_0:SHA_6_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_6_avalon_slave_0_address;              // mm_interconnect_0:SHA_6_avalon_slave_0_address -> SHA_6:address
	wire         mm_interconnect_0_sha_6_avalon_slave_0_write;                // mm_interconnect_0:SHA_6_avalon_slave_0_write -> SHA_6:we
	wire  [31:0] mm_interconnect_0_sha_6_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_6_avalon_slave_0_writedata -> SHA_6:write_data
	wire         mm_interconnect_0_sha_7_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_7_avalon_slave_0_chipselect -> SHA_7:cs
	wire  [31:0] mm_interconnect_0_sha_7_avalon_slave_0_readdata;             // SHA_7:read_data -> mm_interconnect_0:SHA_7_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_7_avalon_slave_0_address;              // mm_interconnect_0:SHA_7_avalon_slave_0_address -> SHA_7:address
	wire         mm_interconnect_0_sha_7_avalon_slave_0_write;                // mm_interconnect_0:SHA_7_avalon_slave_0_write -> SHA_7:we
	wire  [31:0] mm_interconnect_0_sha_7_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_7_avalon_slave_0_writedata -> SHA_7:write_data
	wire         mm_interconnect_0_sha_8_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_8_avalon_slave_0_chipselect -> SHA_8:cs
	wire  [31:0] mm_interconnect_0_sha_8_avalon_slave_0_readdata;             // SHA_8:read_data -> mm_interconnect_0:SHA_8_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_8_avalon_slave_0_address;              // mm_interconnect_0:SHA_8_avalon_slave_0_address -> SHA_8:address
	wire         mm_interconnect_0_sha_8_avalon_slave_0_write;                // mm_interconnect_0:SHA_8_avalon_slave_0_write -> SHA_8:we
	wire  [31:0] mm_interconnect_0_sha_8_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_8_avalon_slave_0_writedata -> SHA_8:write_data
	wire         mm_interconnect_0_sha_9_avalon_slave_0_chipselect;           // mm_interconnect_0:SHA_9_avalon_slave_0_chipselect -> SHA_9:cs
	wire  [31:0] mm_interconnect_0_sha_9_avalon_slave_0_readdata;             // SHA_9:read_data -> mm_interconnect_0:SHA_9_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_sha_9_avalon_slave_0_address;              // mm_interconnect_0:SHA_9_avalon_slave_0_address -> SHA_9:address
	wire         mm_interconnect_0_sha_9_avalon_slave_0_write;                // mm_interconnect_0:SHA_9_avalon_slave_0_write -> SHA_9:we
	wire  [31:0] mm_interconnect_0_sha_9_avalon_slave_0_writedata;            // mm_interconnect_0:SHA_9_avalon_slave_0_writedata -> SHA_9:write_data
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;            // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;              // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_1_s1_address;               // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;            // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                 // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;             // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                 // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire         irq_mapper_receiver10_irq;                                   // jtag_uart_0:av_irq -> irq_mapper:receiver10_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver0_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // SHA_0:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                           // SHA_1:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                    // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                           // SHA_2:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                    // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                           // SHA_3:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver4_irq;                                    // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                           // SHA_4:irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver5_irq;                                    // irq_synchronizer_005:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                           // SHA_5:irq -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver6_irq;                                    // irq_synchronizer_006:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_006_receiver_irq;                           // SHA_6:irq -> irq_synchronizer_006:receiver_irq
	wire         irq_mapper_receiver7_irq;                                    // irq_synchronizer_007:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_007_receiver_irq;                           // SHA_7:irq -> irq_synchronizer_007:receiver_irq
	wire         irq_mapper_receiver8_irq;                                    // irq_synchronizer_008:sender_irq -> irq_mapper:receiver8_irq
	wire   [0:0] irq_synchronizer_008_receiver_irq;                           // SHA_8:irq -> irq_synchronizer_008:receiver_irq
	wire         irq_mapper_receiver9_irq;                                    // irq_synchronizer_009:sender_irq -> irq_mapper:receiver9_irq
	wire   [0:0] irq_synchronizer_009_receiver_irq;                           // SHA_9:irq -> irq_synchronizer_009:receiver_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [SHA_0:reset_n, SHA_1:reset_n, SHA_2:reset_n, SHA_3:reset_n, SHA_4:reset_n, SHA_5:reset_n, SHA_6:reset_n, SHA_7:reset_n, SHA_8:reset_n, SHA_9:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, irq_synchronizer_007:receiver_reset, irq_synchronizer_008:receiver_reset, irq_synchronizer_009:receiver_reset, mm_interconnect_0:SHA_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, irq_synchronizer_008:sender_reset, irq_synchronizer_009:sender_reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, onchip_memory2_1:reset, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]

	sha256 sha_0 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_0_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_0_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_0_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_0_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_0_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_receiver_irq)                      // interrupt_sender.irq
	);

	sha256 sha_1 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_1_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_1_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_1_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_1_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_1_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_001_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_2 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_2_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_2_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_2_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_2_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_2_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_002_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_3 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_3_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_3_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_3_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_3_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_3_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_003_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_4 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_4_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_4_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_4_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_4_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_4_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_004_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_5 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_5_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_5_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_5_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_5_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_5_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_005_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_6 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_6_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_6_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_6_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_6_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_6_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_006_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_7 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_7_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_7_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_7_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_7_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_7_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_007_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_8 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_8_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_8_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_8_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_8_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_8_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_008_receiver_irq)                  // interrupt_sender.irq
	);

	sha256 sha_9 (
		.clk        (pll_0_outclk0_clk),                                 //            clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.we         (mm_interconnect_0_sha_9_avalon_slave_0_write),      //   avalon_slave_0.write
		.address    (mm_interconnect_0_sha_9_avalon_slave_0_address),    //                 .address
		.write_data (mm_interconnect_0_sha_9_avalon_slave_0_writedata),  //                 .writedata
		.read_data  (mm_interconnect_0_sha_9_avalon_slave_0_readdata),   //                 .readdata
		.cs         (mm_interconnect_0_sha_9_avalon_slave_0_chipselect), //                 .chipselect
		.irq        (irq_synchronizer_009_receiver_irq)                  // interrupt_sender.irq
	);

	system_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_clk_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver10_irq)                                    //               irq.irq
	);

	system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sys_clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sys_clk_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	system_onchip_memory2_1 onchip_memory2_1 (
		.clk        (sys_clk_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	system_pll_0 pll_0 (
		.refclk   (sys_clk_clk),       //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   //  locked.export
	);

	system_sdram sdram (
		.clk            (sys_clk_clk),                              //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                              (pll_0_outclk0_clk),                                           //                            pll_0_outclk0.clk
		.system_clk_clk_clk                             (sys_clk_clk),                                                 //                           system_clk_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.SHA_0_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                              //        SHA_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.onchip_memory2_1_s1_address                    (mm_interconnect_0_onchip_memory2_1_s1_address),               //                      onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                      (mm_interconnect_0_onchip_memory2_1_s1_write),                 //                                         .write
		.onchip_memory2_1_s1_readdata                   (mm_interconnect_0_onchip_memory2_1_s1_readdata),              //                                         .readdata
		.onchip_memory2_1_s1_writedata                  (mm_interconnect_0_onchip_memory2_1_s1_writedata),             //                                         .writedata
		.onchip_memory2_1_s1_byteenable                 (mm_interconnect_0_onchip_memory2_1_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_1_s1_chipselect                 (mm_interconnect_0_onchip_memory2_1_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_1_s1_clken                      (mm_interconnect_0_onchip_memory2_1_s1_clken),                 //                                         .clken
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.SHA_0_avalon_slave_0_address                   (mm_interconnect_0_sha_0_avalon_slave_0_address),              //                     SHA_0_avalon_slave_0.address
		.SHA_0_avalon_slave_0_write                     (mm_interconnect_0_sha_0_avalon_slave_0_write),                //                                         .write
		.SHA_0_avalon_slave_0_readdata                  (mm_interconnect_0_sha_0_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_0_avalon_slave_0_writedata                 (mm_interconnect_0_sha_0_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_0_avalon_slave_0_chipselect                (mm_interconnect_0_sha_0_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_1_avalon_slave_0_address                   (mm_interconnect_0_sha_1_avalon_slave_0_address),              //                     SHA_1_avalon_slave_0.address
		.SHA_1_avalon_slave_0_write                     (mm_interconnect_0_sha_1_avalon_slave_0_write),                //                                         .write
		.SHA_1_avalon_slave_0_readdata                  (mm_interconnect_0_sha_1_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_1_avalon_slave_0_writedata                 (mm_interconnect_0_sha_1_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_1_avalon_slave_0_chipselect                (mm_interconnect_0_sha_1_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_2_avalon_slave_0_address                   (mm_interconnect_0_sha_2_avalon_slave_0_address),              //                     SHA_2_avalon_slave_0.address
		.SHA_2_avalon_slave_0_write                     (mm_interconnect_0_sha_2_avalon_slave_0_write),                //                                         .write
		.SHA_2_avalon_slave_0_readdata                  (mm_interconnect_0_sha_2_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_2_avalon_slave_0_writedata                 (mm_interconnect_0_sha_2_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_2_avalon_slave_0_chipselect                (mm_interconnect_0_sha_2_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_3_avalon_slave_0_address                   (mm_interconnect_0_sha_3_avalon_slave_0_address),              //                     SHA_3_avalon_slave_0.address
		.SHA_3_avalon_slave_0_write                     (mm_interconnect_0_sha_3_avalon_slave_0_write),                //                                         .write
		.SHA_3_avalon_slave_0_readdata                  (mm_interconnect_0_sha_3_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_3_avalon_slave_0_writedata                 (mm_interconnect_0_sha_3_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_3_avalon_slave_0_chipselect                (mm_interconnect_0_sha_3_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_4_avalon_slave_0_address                   (mm_interconnect_0_sha_4_avalon_slave_0_address),              //                     SHA_4_avalon_slave_0.address
		.SHA_4_avalon_slave_0_write                     (mm_interconnect_0_sha_4_avalon_slave_0_write),                //                                         .write
		.SHA_4_avalon_slave_0_readdata                  (mm_interconnect_0_sha_4_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_4_avalon_slave_0_writedata                 (mm_interconnect_0_sha_4_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_4_avalon_slave_0_chipselect                (mm_interconnect_0_sha_4_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_5_avalon_slave_0_address                   (mm_interconnect_0_sha_5_avalon_slave_0_address),              //                     SHA_5_avalon_slave_0.address
		.SHA_5_avalon_slave_0_write                     (mm_interconnect_0_sha_5_avalon_slave_0_write),                //                                         .write
		.SHA_5_avalon_slave_0_readdata                  (mm_interconnect_0_sha_5_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_5_avalon_slave_0_writedata                 (mm_interconnect_0_sha_5_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_5_avalon_slave_0_chipselect                (mm_interconnect_0_sha_5_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_6_avalon_slave_0_address                   (mm_interconnect_0_sha_6_avalon_slave_0_address),              //                     SHA_6_avalon_slave_0.address
		.SHA_6_avalon_slave_0_write                     (mm_interconnect_0_sha_6_avalon_slave_0_write),                //                                         .write
		.SHA_6_avalon_slave_0_readdata                  (mm_interconnect_0_sha_6_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_6_avalon_slave_0_writedata                 (mm_interconnect_0_sha_6_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_6_avalon_slave_0_chipselect                (mm_interconnect_0_sha_6_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_7_avalon_slave_0_address                   (mm_interconnect_0_sha_7_avalon_slave_0_address),              //                     SHA_7_avalon_slave_0.address
		.SHA_7_avalon_slave_0_write                     (mm_interconnect_0_sha_7_avalon_slave_0_write),                //                                         .write
		.SHA_7_avalon_slave_0_readdata                  (mm_interconnect_0_sha_7_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_7_avalon_slave_0_writedata                 (mm_interconnect_0_sha_7_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_7_avalon_slave_0_chipselect                (mm_interconnect_0_sha_7_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_8_avalon_slave_0_address                   (mm_interconnect_0_sha_8_avalon_slave_0_address),              //                     SHA_8_avalon_slave_0.address
		.SHA_8_avalon_slave_0_write                     (mm_interconnect_0_sha_8_avalon_slave_0_write),                //                                         .write
		.SHA_8_avalon_slave_0_readdata                  (mm_interconnect_0_sha_8_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_8_avalon_slave_0_writedata                 (mm_interconnect_0_sha_8_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_8_avalon_slave_0_chipselect                (mm_interconnect_0_sha_8_avalon_slave_0_chipselect),           //                                         .chipselect
		.SHA_9_avalon_slave_0_address                   (mm_interconnect_0_sha_9_avalon_slave_0_address),              //                     SHA_9_avalon_slave_0.address
		.SHA_9_avalon_slave_0_write                     (mm_interconnect_0_sha_9_avalon_slave_0_write),                //                                         .write
		.SHA_9_avalon_slave_0_readdata                  (mm_interconnect_0_sha_9_avalon_slave_0_readdata),             //                                         .readdata
		.SHA_9_avalon_slave_0_writedata                 (mm_interconnect_0_sha_9_avalon_slave_0_writedata),            //                                         .writedata
		.SHA_9_avalon_slave_0_chipselect                (mm_interconnect_0_sha_9_avalon_slave_0_chipselect)            //                                         .chipselect
	);

	system_irq_mapper irq_mapper (
		.clk            (sys_clk_clk),                        //        clk.clk
		.reset          (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),           //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),           //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),           //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),           //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),           //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),           //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),           //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),           //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),           //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),           //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),          // receiver10.irq
		.sender_irq     (nios2_gen2_0_irq_irq)                //     sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_007 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_007_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_008 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_008_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver8_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_009 (
		.receiver_clk   (pll_0_outclk0_clk),                  //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_009_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver9_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (sys_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
